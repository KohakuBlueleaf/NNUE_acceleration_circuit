parameter MAX_ROW = 4;
parameter Layer1 = 64;
parameter Layer2 = 16;
parameter Layer3 = 16;