parameter MAX_ROW = 16;
parameter Layer1 = 128;
parameter Layer2 = 16;
parameter Layer3 = 16;