//This project can run in basys3 with MAX_ROW set to 2 
//and use basys3/w2.coe, w3.coe to replace the original w2,w3.coe
parameter MAX_ROW = 2; //use 2 for basys3, 16 for nexys A7
parameter Layer1 = 128;
parameter Layer2 = 16;
parameter Layer3 = 16;