`timescale 1ns/1ps


module VGAController(pclk, reset, hsync, vsync, valid, h_cnt, v_cnt);
    input pclk, reset;
    output hsync, vsync;
	output valid;
    output [9:0]h_cnt, v_cnt;
    
    reg [9:0]pixel_cnt;
    reg [9:0]line_cnt;
    reg hsync_i,vsync_i;
	wire hsync_default, vsync_default;
    wire [9:0] HD, HF, HS, HB, HT, VD, VF, VS, VB, VT;
	
    assign HD = 640;
    assign HF = 16;
    assign HS = 96;
    assign HB = 48;
    assign HT = 800; 
    assign VD = 480;
    assign VF = 10;
    assign VS = 2;
    assign VB = 33;
    assign VT = 525;
    assign hsync_default = 1'b1;
    assign vsync_default = 1'b1;
    
    always@(posedge pclk)
        if(reset)
            pixel_cnt <= 0;
        else if(pixel_cnt < (HT - 1))
            pixel_cnt <= pixel_cnt + 1;
        else
            pixel_cnt <= 0;

    always@(posedge pclk)
        if(reset)
            hsync_i <= hsync_default;
        else if((pixel_cnt >= (HD + HF - 1))&&(pixel_cnt < (HD + HF + HS - 1)))
                hsync_i <= ~hsync_default;
            else
                hsync_i <= hsync_default; 
    
    always@(posedge pclk)
        if(reset)
            line_cnt <= 0;
        else if(pixel_cnt == (HT -1))
            if(line_cnt < (VT - 1))
                line_cnt <= line_cnt + 1;
            else
                line_cnt <= 0;
        else
            line_cnt <= line_cnt;
    
    
    always@(posedge pclk)
        if(reset)
            vsync_i <= vsync_default; 
        else if((line_cnt >= (VD + VF - 1))&&(line_cnt < (VD + VF + VS - 1)))
            vsync_i <= ~vsync_default;
        else
            vsync_i <= vsync_default; 

    assign hsync = hsync_i;
    assign vsync = vsync_i;
    assign valid = ((pixel_cnt < HD) && (line_cnt < VD));

    assign h_cnt = (pixel_cnt < HD)? pixel_cnt : 10'd0;//639
    assign v_cnt = (line_cnt < VD)? line_cnt : 10'd0;//479
endmodule


module DisplayVGA(
    input clk, rst, 
    input player,               // Which player takes control (matained by Status)
    input [1:0] game_status,    // Game status generated by Status
    input [7:0] addr0, addr1,   // Address generated by Input
    input [0:241] board,        // Board maintained by Status
    input [0:120] win_board,    // Win chesses position maintained by Status
    input [15:0] score,         // The score generated by NNUE
    output [3:0] vgaRed, vgaBlue, vgaGreen,
    output [9:0] shift,
    output hsync, vsync
);  
    // RGB color assignment
    parameter BG = 12'hddd;
    parameter BOARD = 12'hfcd;
    parameter GRID = 12'h8a8;
    parameter SCORE = 12'h659;
    parameter BLACK = 12'h000;
    parameter WHITE = 12'hFFF;
    parameter PURPLE = 12'h409;
    parameter RED   = 12'hD22;
    parameter GRAY  = 12'h555;
    parameter BLUE  = 12'h58A;

    reg [11:0] usedcolor, next_usedcolor;
    assign {vgaRed, vgaGreen, vgaBlue} = (valid) ? usedcolor : BLACK;

    always @(posedge clk) begin
        if (rst) begin
            usedcolor <= BLACK;
        end else begin
            usedcolor <= next_usedcolor;
        end
    end

    // vga controller
    wire valid;
    wire [9:0] h_cnt, v_cnt;
    VGAController VC0 (
        .pclk(clk),
        .reset(rst),
        .hsync(hsync),
        .vsync(vsync),
        .valid(valid),
        .h_cnt(h_cnt),
        .v_cnt(v_cnt)
    );    

    // Chessboard infomation
    parameter CHESS_RADIUS = 10;
    parameter PADDING = 4;
    parameter BLOCK_WIDTH = 2 * CHESS_RADIUS + 2 * PADDING;
    parameter LINE_WIDTH = 4;
    parameter BOARD_WIDTH = 11 * (BLOCK_WIDTH) + 12 * LINE_WIDTH;
    parameter BOARD_H = 140;
    parameter BOARD_V = 40;
    parameter SCORE_H = BOARD_H;
    parameter SCORE_V = BOARD_V + BOARD_WIDTH + 20;
    parameter SCORE_H_LEN = BOARD_WIDTH;
    parameter SCORE_V_LEN = 30;
    parameter SCORE_MAX = 6000;

    // Usedcolor update
    wire [3:0] block_v, block_h, chess_h, chess_v;
    wire [7:0] blockaddr0, blockaddr1;
    wire [15:0] blockmid_v_cnt, blockmid_h_cnt, v_diff, h_diff;
    wire [15:0] abs_score, clipped, ratio;
    wire [9:0] shift; // calculate the shift from the mid point of score.
    wire [9:0] score_div_pt; // h_cnt <= score_div_pt will represent the score for white, vise versa.
    wire in_chessboard, in_line, draw_rec, in_chess, in_score, in_score_mid;

    assign chess_v          = addr0 / 11;
    assign chess_h          = addr0 % 11;
    assign block_v          = (v_cnt - BOARD_V) / (BLOCK_WIDTH + LINE_WIDTH); // Index of v of current block.
    assign block_h          = (h_cnt - BOARD_H) / (BLOCK_WIDTH + LINE_WIDTH); // Index of h of current block.
    assign blockaddr0       = block_v * 11 + block_h;
    assign blockaddr1       = blockaddr0 + 8'd121;
    assign blockmid_v_cnt   = BOARD_V + block_v * (BLOCK_WIDTH + LINE_WIDTH) + LINE_WIDTH + BLOCK_WIDTH / 2; // Pixel of v of midpoint of current block
    assign blockmid_h_cnt   = BOARD_H + block_h * (BLOCK_WIDTH + LINE_WIDTH) + LINE_WIDTH + BLOCK_WIDTH / 2; // Pixel of h of midpoint of current block
    assign v_diff           = (blockmid_v_cnt > v_cnt) ? blockmid_v_cnt - v_cnt : v_cnt - blockmid_v_cnt;
    assign h_diff           = (blockmid_h_cnt > h_cnt) ? blockmid_h_cnt - h_cnt : h_cnt - blockmid_h_cnt;
    assign in_chessboard    = (h_cnt >= BOARD_H && h_cnt < BOARD_H + BOARD_WIDTH) && (v_cnt >= BOARD_V && v_cnt < BOARD_V + BOARD_WIDTH); // Whether the pixel is in the chessboard
    assign in_line          = ((h_cnt - BOARD_H) % (BLOCK_WIDTH + LINE_WIDTH) < LINE_WIDTH) || ((v_cnt - BOARD_V) % (BLOCK_WIDTH + LINE_WIDTH) < LINE_WIDTH); // Whether the pixel is in the line
    assign draw_rec         = (game_status == 0) && in_line && (
                                (block_v == chess_v && block_h == chess_h) ||
                                (block_v == chess_v + 1 && block_h == chess_h && v_cnt < blockmid_v_cnt - BLOCK_WIDTH / 2) ||
                                (block_v == chess_v && block_h == chess_h + 1 && h_cnt < blockmid_h_cnt - BLOCK_WIDTH / 2) ||
                                (block_v == chess_v + 1 && block_h == chess_h + 1 && h_cnt < blockmid_h_cnt - BLOCK_WIDTH / 2 && v_cnt < blockmid_v_cnt - BLOCK_WIDTH / 2)
                            );
    assign in_chess         = (h_diff * h_diff + v_diff * v_diff < CHESS_RADIUS * CHESS_RADIUS);
    assign in_score         = (SCORE_H <= h_cnt && h_cnt <= SCORE_H + SCORE_H_LEN) && (SCORE_V <= v_cnt && v_cnt <= SCORE_V + SCORE_V_LEN);
    assign in_score_mid     = (SCORE_H + PADDING <= h_cnt && h_cnt + PADDING <= SCORE_H + SCORE_H_LEN) && (SCORE_V + PADDING <= v_cnt && v_cnt + PADDING <= SCORE_V + SCORE_V_LEN);
    assign abs_score        = (score[15]) ? ~(score - 1) : score;
    assign clipped          = (abs_score > SCORE_MAX) ? SCORE_MAX : abs_score;
    assign ratio            = SCORE_MAX * 2 / SCORE_H_LEN;
    assign shift            = (clipped / ratio > SCORE_H_LEN / 2) ? SCORE_H_LEN / 2 : clipped / ratio; // abs_score
    assign score_div_pt     = (game_status == 2'b01) ? SCORE_H + SCORE_H_LEN - PADDING :(
                                (game_status == 2'b10) ? SCORE_H :(
                                ~(score[15] ^ player) ? SCORE_H + SCORE_H_LEN / 2 + shift : SCORE_H + SCORE_H_LEN / 2 - shift
                                )
                            ); 

    // next_usedcolor assignment
    always @(*) begin
        if (in_chessboard) begin
            if (~in_line) begin
                if (in_chess) begin 
                    if (game_status) begin
                        case({board[blockaddr0], board[blockaddr1], win_board[blockaddr0]})
                            3'b011: next_usedcolor = BLACK;
                            3'b101: next_usedcolor = WHITE;
                            default: next_usedcolor = BOARD;
                        endcase
                    end else begin
                        case({board[blockaddr0], board[blockaddr1]}) // First hand will be white
                            2'b01: next_usedcolor = BLACK;
                            2'b10: next_usedcolor = WHITE;
                            default: next_usedcolor = BOARD;
                        endcase       
                    end             
                end else
                    next_usedcolor = BOARD;
            end else begin
                next_usedcolor = draw_rec ? (player ? BLACK : WHITE) : GRID;
            end
        end else if (in_score) begin
            if (in_score_mid) begin
                next_usedcolor = (h_cnt <= score_div_pt) ? WHITE : BLACK;
            end else begin
                next_usedcolor = SCORE;
            end
        end else begin
            next_usedcolor = BG;
        end
    end
endmodule